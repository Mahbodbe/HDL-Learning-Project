library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Top_indirect is
    Port ( unlock, cunlock, reset, vcc_1, s_i : in  STD_LOGIC;
           clk, clk_d : in  STD_LOGIC;
           y : out  STD_LOGIC);
end Top_indirect;

architecture Behavioral of Top_indirect is

component counter is
	generic
	(
	   num :integer
	);
    Port ( clk : in  STD_LOGIC;
           reset : in  STD_LOGIC;
           Outc : out  STD_LOGIC_VECTOR (num -1 downto 0));
end component;

component Comparator16 is
    Port ( Ac, Bc : in  STD_LOGIC_VECTOR (15 downto 0);
           Oc : out  STD_LOGIC);
end component;

component JKFF is
    Port (
        K, J   : in  STD_LOGIC;
        clk    : in  STD_LOGIC;
        reset  : in  STD_LOGIC;
        Ojk    : out STD_LOGIC
    );
end component;

component Sync_D_FlipFlop is
    Port ( D : in  STD_LOGIC;
           clk : in  STD_LOGIC;
           reset : in  STD_LOGIC;
           Q : out  STD_LOGIC);
end component;


component Mux2x1 is
    Port ( Am2 : in  STD_LOGIC_VECTOR (1 downto 0);
           Om2 : out  STD_LOGIC;
           Sm2 : in  STD_LOGIC);
end component;

component Mux8x1 is
    Port ( Am : in  STD_LOGIC_VECTOR (7 downto 0);
           Om : out  STD_LOGIC;
           Sm : in  STD_LOGIC_VECTOR (2 downto 0));
end component;

component SIPO_parametric is
	generic 
	(
		number:integer
	);
    Port ( si : in  STD_LOGIC;
           clk : in  STD_LOGIC;
           res : in  STD_LOGIC;
           Osipo : out  STD_LOGIC_VECTOR (number-1 downto 0));
end component;


signal unlock_b, cunlock_b, reset_b, jclk, js, k, M1, M2, b1, DO : STD_LOGIC :='0';
signal q : STD_LOGIC_VECTOR(31 downto 0) := (others => '0');
signal x : STD_LOGIC_VECTOR(2 downto 0) := (others => '0');
signal O8 : STD_LOGIC_VECTOR(7 downto 0) := (others => '0');
signal CA, CB : STD_LOGIC_VECTOR(15 downto 0) := (others => '0');
signal reset_u3, clk_u4, reset_u5 : STD_LOGIC := '0';



begin

unlock_b <= not unlock;
cunlock_b <= not cunlock;
reset_b <= not reset; 
reset_u3 <= unlock_b or reset_b;
clk_u4 <= b1 and (not DO);
reset_u5 <= reset_b or jclk;

u1:counter generic map ( num => 32) port map (clk => clk, reset => reset_b, Outc=> q );
u2:Comparator16 port map ( Ac => CA, Bc => CB, Oc => jclk);
u3: JKFF port map (K => '1', J => js, clk => jclk, Ojk => k, reset => reset_u3);
u4: counter generic map (num => 3) port map (clk => clk_u4, reset => reset_b, Outc => x);
u5: counter generic map (num => 16) port map (clk => M1, reset => reset_u5, Outc => CA);
u6:Sync_D_FlipFlop port map(D => b1, Q => DO, reset => reset_b, clk => q(11));
u7:Mux2x1 port map(Am2(0) => '1', Am2(1) => '0', Sm2 => cunlock_b, Om2 => js);
u8:Mux2x1 port map(Am2(0) => M2, Am2(1) => '0', Sm2 => k, Om2=> M1);
u9:Mux8x1 port map(Am(0) => q(31), Am(1) => q(27), Am(2) => q(23), Am(3) => q(19), Am(4) => q(15), Am(5) => q(11), Am(6) => q(7), Am(7) => q(3), Om => M2, Sm=> x);
u10:SIPO_parametric generic map (number => 16) port map(si => s_i, clk => clk_d, res => reset_b, Osipo => CB);
u11:SIPO_parametric generic map (number => 8) port map(si => vcc_1, clk => q(11), res => reset_b, Osipo => O8);
b1 <= O8(0) and O8(1) and O8(2) and O8(3) and O8(4) and O8(5) and O8(6) and O8(7);
y <= k;


end Behavioral;

