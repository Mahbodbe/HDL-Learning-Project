`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    08:17:34 05/12/2025 
// Design Name: 
// Module Name:    FB_Async_sync_D_FF 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module FB_Async_sync_D_FF(
    input [3:0] D_FB,
    input reset_fb,
    input set_fb,
    input clk,
    output [3:0] Q_FB
    );


endmodule
